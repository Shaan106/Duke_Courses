module divider_superfast(
    data_operandA, data_operandB, 
    clock, 
    data_result, data_exception, data_resultRDY);

    input [31:0] data_operandA, data_operandB;
    input clock;

    output [63:0] data_result;
    output data_exception, data_resultRDY;

    //COUNTER COUNTER
    

endmodule